// onchip_ram_256b.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module onchip_ram_256b (
		input  wire         clk_clk,                        //              clk.clk
		output wire         host_bridge_1_s0_waitrequest,   // host_bridge_1_s0.waitrequest
		output wire [255:0] host_bridge_1_s0_readdata,      //                 .readdata
		output wire         host_bridge_1_s0_readdatavalid, //                 .readdatavalid
		input  wire [0:0]   host_bridge_1_s0_burstcount,    //                 .burstcount
		input  wire [255:0] host_bridge_1_s0_writedata,     //                 .writedata
		input  wire [22:0]  host_bridge_1_s0_address,       //                 .address
		input  wire         host_bridge_1_s0_write,         //                 .write
		input  wire         host_bridge_1_s0_read,          //                 .read
		input  wire [31:0]  host_bridge_1_s0_byteenable,    //                 .byteenable
		input  wire         host_bridge_1_s0_debugaccess,   //                 .debugaccess
		output wire         kernel_bridge_s0_waitrequest,   // kernel_bridge_s0.waitrequest
		output wire [255:0] kernel_bridge_s0_readdata,      //                 .readdata
		output wire         kernel_bridge_s0_readdatavalid, //                 .readdatavalid
		input  wire [4:0]   kernel_bridge_s0_burstcount,    //                 .burstcount
		input  wire [255:0] kernel_bridge_s0_writedata,     //                 .writedata
		input  wire [22:0]  kernel_bridge_s0_address,       //                 .address
		input  wire         kernel_bridge_s0_write,         //                 .write
		input  wire         kernel_bridge_s0_read,          //                 .read
		input  wire [31:0]  kernel_bridge_s0_byteenable,    //                 .byteenable
		input  wire         kernel_bridge_s0_debugaccess,   //                 .debugaccess
		input  wire         reset_reset_n                   //            reset.reset_n
	);

	wire          host_bridge_1_m0_waitrequest;                     // mm_interconnect_0:host_bridge_1_m0_waitrequest -> host_bridge_1:m0_waitrequest
	wire  [255:0] host_bridge_1_m0_readdata;                        // mm_interconnect_0:host_bridge_1_m0_readdata -> host_bridge_1:m0_readdata
	wire          host_bridge_1_m0_debugaccess;                     // host_bridge_1:m0_debugaccess -> mm_interconnect_0:host_bridge_1_m0_debugaccess
	wire   [22:0] host_bridge_1_m0_address;                         // host_bridge_1:m0_address -> mm_interconnect_0:host_bridge_1_m0_address
	wire          host_bridge_1_m0_read;                            // host_bridge_1:m0_read -> mm_interconnect_0:host_bridge_1_m0_read
	wire   [31:0] host_bridge_1_m0_byteenable;                      // host_bridge_1:m0_byteenable -> mm_interconnect_0:host_bridge_1_m0_byteenable
	wire          host_bridge_1_m0_readdatavalid;                   // mm_interconnect_0:host_bridge_1_m0_readdatavalid -> host_bridge_1:m0_readdatavalid
	wire  [255:0] host_bridge_1_m0_writedata;                       // host_bridge_1:m0_writedata -> mm_interconnect_0:host_bridge_1_m0_writedata
	wire          host_bridge_1_m0_write;                           // host_bridge_1:m0_write -> mm_interconnect_0:host_bridge_1_m0_write
	wire    [0:0] host_bridge_1_m0_burstcount;                      // host_bridge_1:m0_burstcount -> mm_interconnect_0:host_bridge_1_m0_burstcount
	wire          kernel_bridge_m0_waitrequest;                     // mm_interconnect_0:kernel_bridge_m0_waitrequest -> kernel_bridge:m0_waitrequest
	wire  [255:0] kernel_bridge_m0_readdata;                        // mm_interconnect_0:kernel_bridge_m0_readdata -> kernel_bridge:m0_readdata
	wire          kernel_bridge_m0_debugaccess;                     // kernel_bridge:m0_debugaccess -> mm_interconnect_0:kernel_bridge_m0_debugaccess
	wire   [22:0] kernel_bridge_m0_address;                         // kernel_bridge:m0_address -> mm_interconnect_0:kernel_bridge_m0_address
	wire          kernel_bridge_m0_read;                            // kernel_bridge:m0_read -> mm_interconnect_0:kernel_bridge_m0_read
	wire   [31:0] kernel_bridge_m0_byteenable;                      // kernel_bridge:m0_byteenable -> mm_interconnect_0:kernel_bridge_m0_byteenable
	wire          kernel_bridge_m0_readdatavalid;                   // mm_interconnect_0:kernel_bridge_m0_readdatavalid -> kernel_bridge:m0_readdatavalid
	wire  [255:0] kernel_bridge_m0_writedata;                       // kernel_bridge:m0_writedata -> mm_interconnect_0:kernel_bridge_m0_writedata
	wire          kernel_bridge_m0_write;                           // kernel_bridge:m0_write -> mm_interconnect_0:kernel_bridge_m0_write
	wire    [4:0] kernel_bridge_m0_burstcount;                      // kernel_bridge:m0_burstcount -> mm_interconnect_0:kernel_bridge_m0_burstcount
	wire          mm_interconnect_0_onchip_memory2_0_s1_chipselect; // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [255:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;   // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [17:0] mm_interconnect_0_onchip_memory2_0_s1_address;    // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [31:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable; // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire          mm_interconnect_0_onchip_memory2_0_s1_write;      // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [255:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;  // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire          mm_interconnect_0_onchip_memory2_0_s1_clken;      // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire          rst_controller_reset_out_reset;                   // rst_controller:reset_out -> [host_bridge_1:reset, kernel_bridge:reset, mm_interconnect_0:host_bridge_1_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset]

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (256),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (23),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) host_bridge_1 (
		.clk              (clk_clk),                        //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (host_bridge_1_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (host_bridge_1_s0_readdata),      //      .readdata
		.s0_readdatavalid (host_bridge_1_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (host_bridge_1_s0_burstcount),    //      .burstcount
		.s0_writedata     (host_bridge_1_s0_writedata),     //      .writedata
		.s0_address       (host_bridge_1_s0_address),       //      .address
		.s0_write         (host_bridge_1_s0_write),         //      .write
		.s0_read          (host_bridge_1_s0_read),          //      .read
		.s0_byteenable    (host_bridge_1_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (host_bridge_1_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (host_bridge_1_m0_waitrequest),   //    m0.waitrequest
		.m0_readdata      (host_bridge_1_m0_readdata),      //      .readdata
		.m0_readdatavalid (host_bridge_1_m0_readdatavalid), //      .readdatavalid
		.m0_burstcount    (host_bridge_1_m0_burstcount),    //      .burstcount
		.m0_writedata     (host_bridge_1_m0_writedata),     //      .writedata
		.m0_address       (host_bridge_1_m0_address),       //      .address
		.m0_write         (host_bridge_1_m0_write),         //      .write
		.m0_read          (host_bridge_1_m0_read),          //      .read
		.m0_byteenable    (host_bridge_1_m0_byteenable),    //      .byteenable
		.m0_debugaccess   (host_bridge_1_m0_debugaccess),   //      .debugaccess
		.s0_response      (),                               // (terminated)
		.m0_response      (2'b00)                           // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (256),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (23),
		.BURSTCOUNT_WIDTH  (5),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) kernel_bridge (
		.clk              (clk_clk),                        //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (kernel_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (kernel_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (kernel_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (kernel_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (kernel_bridge_s0_writedata),     //      .writedata
		.s0_address       (kernel_bridge_s0_address),       //      .address
		.s0_write         (kernel_bridge_s0_write),         //      .write
		.s0_read          (kernel_bridge_s0_read),          //      .read
		.s0_byteenable    (kernel_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (kernel_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (kernel_bridge_m0_waitrequest),   //    m0.waitrequest
		.m0_readdata      (kernel_bridge_m0_readdata),      //      .readdata
		.m0_readdatavalid (kernel_bridge_m0_readdatavalid), //      .readdatavalid
		.m0_burstcount    (kernel_bridge_m0_burstcount),    //      .burstcount
		.m0_writedata     (kernel_bridge_m0_writedata),     //      .writedata
		.m0_address       (kernel_bridge_m0_address),       //      .address
		.m0_write         (kernel_bridge_m0_write),         //      .write
		.m0_read          (kernel_bridge_m0_read),          //      .read
		.m0_byteenable    (kernel_bridge_m0_byteenable),    //      .byteenable
		.m0_debugaccess   (kernel_bridge_m0_debugaccess),   //      .debugaccess
		.s0_response      (),                               // (terminated)
		.m0_response      (2'b00)                           // (terminated)
	);

	onchip_ram_256b_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (1'b0)                                              // (terminated)
	);

	onchip_ram_256b_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                   (clk_clk),                                          //                                 clk_0_clk.clk
		.host_bridge_1_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // host_bridge_1_reset_reset_bridge_in_reset.reset
		.host_bridge_1_m0_address                        (host_bridge_1_m0_address),                         //                          host_bridge_1_m0.address
		.host_bridge_1_m0_waitrequest                    (host_bridge_1_m0_waitrequest),                     //                                          .waitrequest
		.host_bridge_1_m0_burstcount                     (host_bridge_1_m0_burstcount),                      //                                          .burstcount
		.host_bridge_1_m0_byteenable                     (host_bridge_1_m0_byteenable),                      //                                          .byteenable
		.host_bridge_1_m0_read                           (host_bridge_1_m0_read),                            //                                          .read
		.host_bridge_1_m0_readdata                       (host_bridge_1_m0_readdata),                        //                                          .readdata
		.host_bridge_1_m0_readdatavalid                  (host_bridge_1_m0_readdatavalid),                   //                                          .readdatavalid
		.host_bridge_1_m0_write                          (host_bridge_1_m0_write),                           //                                          .write
		.host_bridge_1_m0_writedata                      (host_bridge_1_m0_writedata),                       //                                          .writedata
		.host_bridge_1_m0_debugaccess                    (host_bridge_1_m0_debugaccess),                     //                                          .debugaccess
		.kernel_bridge_m0_address                        (kernel_bridge_m0_address),                         //                          kernel_bridge_m0.address
		.kernel_bridge_m0_waitrequest                    (kernel_bridge_m0_waitrequest),                     //                                          .waitrequest
		.kernel_bridge_m0_burstcount                     (kernel_bridge_m0_burstcount),                      //                                          .burstcount
		.kernel_bridge_m0_byteenable                     (kernel_bridge_m0_byteenable),                      //                                          .byteenable
		.kernel_bridge_m0_read                           (kernel_bridge_m0_read),                            //                                          .read
		.kernel_bridge_m0_readdata                       (kernel_bridge_m0_readdata),                        //                                          .readdata
		.kernel_bridge_m0_readdatavalid                  (kernel_bridge_m0_readdatavalid),                   //                                          .readdatavalid
		.kernel_bridge_m0_write                          (kernel_bridge_m0_write),                           //                                          .write
		.kernel_bridge_m0_writedata                      (kernel_bridge_m0_writedata),                       //                                          .writedata
		.kernel_bridge_m0_debugaccess                    (kernel_bridge_m0_debugaccess),                     //                                          .debugaccess
		.onchip_memory2_0_s1_address                     (mm_interconnect_0_onchip_memory2_0_s1_address),    //                       onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                       (mm_interconnect_0_onchip_memory2_0_s1_write),      //                                          .write
		.onchip_memory2_0_s1_readdata                    (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //                                          .readdata
		.onchip_memory2_0_s1_writedata                   (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //                                          .writedata
		.onchip_memory2_0_s1_byteenable                  (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //                                          .byteenable
		.onchip_memory2_0_s1_chipselect                  (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //                                          .chipselect
		.onchip_memory2_0_s1_clken                       (mm_interconnect_0_onchip_memory2_0_s1_clken)       //                                          .clken
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
